//-----------------------------------------------------------------------------
// This is used for testing
//-----------------------------------------------------------------------------
